// megafunction wizard: %LPM_LATCH%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_latch 

// ============================================================
// File Name: lpm_latch2.v
// Megafunction Name(s):
// 			lpm_latch
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 222 10/21/2009 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2009 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module lpm_latch2 (
	data,
	gate,
	q);

	input	  data;
	input	  gate;
	output	  q;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: aclr NUMERIC "0"
// Retrieval info: PRIVATE: aset NUMERIC "0"
// Retrieval info: PRIVATE: nBit NUMERIC "1"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_LATCH"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "1"
// Retrieval info: USED_PORT: data 0 0 0 0 INPUT NODEFVAL data
// Retrieval info: USED_PORT: gate 0 0 0 0 INPUT NODEFVAL gate
// Retrieval info: USED_PORT: q 0 0 0 0 OUTPUT NODEFVAL q
// Retrieval info: CONNECT: @data 0 0 1 0 data 0 0 0 0
// Retrieval info: CONNECT: q 0 0 0 0 @q 0 0 1 0
// Retrieval info: CONNECT: @gate 0 0 0 0 gate 0 0 0 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch2.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch2.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch2.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch2.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch2_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_latch2_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
