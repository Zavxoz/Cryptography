// megafunction wizard: %LPM_CONSTANT%VBB%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_constant 

// ============================================================
// File Name: lpm_constantpaddleng.v
// Megafunction Name(s):
// 			lpm_constant
//
// Simulation Library Files(s):
// 			
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 222 10/21/2009 SJ Full Version
// ************************************************************

//Copyright (C) 1991-2009 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.

module lpm_constantpaddleng (
	result)/* synthesis synthesis_clearbox = 1 */;

	output	[255:0]  result;

endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: JTAG_ENABLED NUMERIC "0"
// Retrieval info: PRIVATE: JTAG_ID STRING "NONE"
// Retrieval info: PRIVATE: Radix NUMERIC "16"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: PRIVATE: Value NUMERIC "640"
// Retrieval info: PRIVATE: nBit NUMERIC "256"
// Retrieval info: CONSTANT: LPM_CVALUE NUMERIC "640"
// Retrieval info: CONSTANT: LPM_HINT STRING "ENABLE_RUNTIME_MOD=NO"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_CONSTANT"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "256"
// Retrieval info: USED_PORT: result 0 0 256 0 OUTPUT NODEFVAL result[255..0]
// Retrieval info: CONNECT: result 0 0 256 0 @result 0 0 256 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_constantpaddleng.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_constantpaddleng.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_constantpaddleng.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_constantpaddleng.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_constantpaddleng_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_constantpaddleng_bb.v TRUE
