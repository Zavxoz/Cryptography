// megafunction wizard: %LPM_MUX%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: lpm_mux 

// ============================================================
// File Name: lpm_mux641.v
// Megafunction Name(s):
// 			lpm_mux
//
// Simulation Library Files(s):
// 			lpm
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 9.1 Build 222 10/21/2009 SJ Full Version
// ************************************************************


//Copyright (C) 1991-2009 Altera Corporation
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, Altera MegaCore Function License 
//Agreement, or other applicable license agreement, including, 
//without limitation, that your use is for the sole purpose of 
//programming logic devices manufactured by Altera and sold by 
//Altera or its authorized distributors.  Please refer to the 
//applicable agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module lpm_mux641 (
	data0,
	data1,
	data10,
	data11,
	data12,
	data13,
	data14,
	data15,
	data16,
	data17,
	data18,
	data19,
	data2,
	data20,
	data21,
	data22,
	data23,
	data24,
	data25,
	data26,
	data27,
	data28,
	data29,
	data3,
	data30,
	data31,
	data32,
	data33,
	data34,
	data35,
	data36,
	data37,
	data38,
	data39,
	data4,
	data40,
	data41,
	data42,
	data43,
	data44,
	data45,
	data46,
	data47,
	data48,
	data49,
	data5,
	data50,
	data51,
	data52,
	data53,
	data54,
	data55,
	data56,
	data57,
	data58,
	data59,
	data6,
	data60,
	data61,
	data62,
	data63,
	data7,
	data8,
	data9,
	sel,
	result);

	input	  data0;
	input	  data1;
	input	  data10;
	input	  data11;
	input	  data12;
	input	  data13;
	input	  data14;
	input	  data15;
	input	  data16;
	input	  data17;
	input	  data18;
	input	  data19;
	input	  data2;
	input	  data20;
	input	  data21;
	input	  data22;
	input	  data23;
	input	  data24;
	input	  data25;
	input	  data26;
	input	  data27;
	input	  data28;
	input	  data29;
	input	  data3;
	input	  data30;
	input	  data31;
	input	  data32;
	input	  data33;
	input	  data34;
	input	  data35;
	input	  data36;
	input	  data37;
	input	  data38;
	input	  data39;
	input	  data4;
	input	  data40;
	input	  data41;
	input	  data42;
	input	  data43;
	input	  data44;
	input	  data45;
	input	  data46;
	input	  data47;
	input	  data48;
	input	  data49;
	input	  data5;
	input	  data50;
	input	  data51;
	input	  data52;
	input	  data53;
	input	  data54;
	input	  data55;
	input	  data56;
	input	  data57;
	input	  data58;
	input	  data59;
	input	  data6;
	input	  data60;
	input	  data61;
	input	  data62;
	input	  data63;
	input	  data7;
	input	  data8;
	input	  data9;
	input	[5:0]  sel;
	output	  result;

	wire [0:0] sub_wire0;
	wire  sub_wire66 = data63;
	wire  sub_wire65 = data61;
	wire  sub_wire64 = data60;
	wire  sub_wire63 = data59;
	wire  sub_wire62 = data58;
	wire  sub_wire61 = data57;
	wire  sub_wire60 = data56;
	wire  sub_wire59 = data55;
	wire  sub_wire58 = data54;
	wire  sub_wire57 = data53;
	wire  sub_wire56 = data52;
	wire  sub_wire55 = data51;
	wire  sub_wire54 = data50;
	wire  sub_wire53 = data49;
	wire  sub_wire52 = data48;
	wire  sub_wire51 = data47;
	wire  sub_wire50 = data46;
	wire  sub_wire49 = data45;
	wire  sub_wire48 = data44;
	wire  sub_wire47 = data43;
	wire  sub_wire46 = data42;
	wire  sub_wire45 = data41;
	wire  sub_wire44 = data40;
	wire  sub_wire43 = data39;
	wire  sub_wire42 = data38;
	wire  sub_wire41 = data37;
	wire  sub_wire40 = data36;
	wire  sub_wire39 = data35;
	wire  sub_wire38 = data34;
	wire  sub_wire37 = data33;
	wire  sub_wire36 = data32;
	wire  sub_wire35 = data31;
	wire  sub_wire34 = data30;
	wire  sub_wire33 = data29;
	wire  sub_wire32 = data28;
	wire  sub_wire31 = data27;
	wire  sub_wire30 = data26;
	wire  sub_wire29 = data25;
	wire  sub_wire28 = data24;
	wire  sub_wire27 = data23;
	wire  sub_wire26 = data22;
	wire  sub_wire25 = data21;
	wire  sub_wire24 = data20;
	wire  sub_wire23 = data19;
	wire  sub_wire22 = data18;
	wire  sub_wire21 = data17;
	wire  sub_wire20 = data16;
	wire  sub_wire19 = data15;
	wire  sub_wire18 = data14;
	wire  sub_wire17 = data13;
	wire  sub_wire16 = data12;
	wire  sub_wire15 = data11;
	wire  sub_wire14 = data10;
	wire  sub_wire13 = data9;
	wire  sub_wire12 = data8;
	wire  sub_wire11 = data7;
	wire  sub_wire10 = data6;
	wire  sub_wire9 = data5;
	wire  sub_wire8 = data4;
	wire  sub_wire7 = data3;
	wire  sub_wire6 = data2;
	wire  sub_wire5 = data1;
	wire  sub_wire4 = data0;
	wire [0:0] sub_wire1 = sub_wire0[0:0];
	wire  result = sub_wire1;
	wire  sub_wire2 = data62;
	wire [63:0] sub_wire3 = {sub_wire66, sub_wire2, sub_wire65, sub_wire64, sub_wire63, sub_wire62, sub_wire61, sub_wire60, sub_wire59, sub_wire58, sub_wire57, sub_wire56, sub_wire55, sub_wire54, sub_wire53, sub_wire52, sub_wire51, sub_wire50, sub_wire49, sub_wire48, sub_wire47, sub_wire46, sub_wire45, sub_wire44, sub_wire43, sub_wire42, sub_wire41, sub_wire40, sub_wire39, sub_wire38, sub_wire37, sub_wire36, sub_wire35, sub_wire34, sub_wire33, sub_wire32, sub_wire31, sub_wire30, sub_wire29, sub_wire28, sub_wire27, sub_wire26, sub_wire25, sub_wire24, sub_wire23, sub_wire22, sub_wire21, sub_wire20, sub_wire19, sub_wire18, sub_wire17, sub_wire16, sub_wire15, sub_wire14, sub_wire13, sub_wire12, sub_wire11, sub_wire10, sub_wire9, sub_wire8, sub_wire7, sub_wire6, sub_wire5, sub_wire4};

	lpm_mux	lpm_mux_component (
				.sel (sel),
				.data (sub_wire3),
				.result (sub_wire0)
				// synopsys translate_off
				,
				.aclr (),
				.clken (),
				.clock ()
				// synopsys translate_on
				);
	defparam
		lpm_mux_component.lpm_size = 64,
		lpm_mux_component.lpm_type = "LPM_MUX",
		lpm_mux_component.lpm_width = 1,
		lpm_mux_component.lpm_widths = 6;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone II"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: CONSTANT: LPM_SIZE NUMERIC "64"
// Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
// Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "1"
// Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "6"
// Retrieval info: USED_PORT: data0 0 0 0 0 INPUT NODEFVAL data0
// Retrieval info: USED_PORT: data1 0 0 0 0 INPUT NODEFVAL data1
// Retrieval info: USED_PORT: data10 0 0 0 0 INPUT NODEFVAL data10
// Retrieval info: USED_PORT: data11 0 0 0 0 INPUT NODEFVAL data11
// Retrieval info: USED_PORT: data12 0 0 0 0 INPUT NODEFVAL data12
// Retrieval info: USED_PORT: data13 0 0 0 0 INPUT NODEFVAL data13
// Retrieval info: USED_PORT: data14 0 0 0 0 INPUT NODEFVAL data14
// Retrieval info: USED_PORT: data15 0 0 0 0 INPUT NODEFVAL data15
// Retrieval info: USED_PORT: data16 0 0 0 0 INPUT NODEFVAL data16
// Retrieval info: USED_PORT: data17 0 0 0 0 INPUT NODEFVAL data17
// Retrieval info: USED_PORT: data18 0 0 0 0 INPUT NODEFVAL data18
// Retrieval info: USED_PORT: data19 0 0 0 0 INPUT NODEFVAL data19
// Retrieval info: USED_PORT: data2 0 0 0 0 INPUT NODEFVAL data2
// Retrieval info: USED_PORT: data20 0 0 0 0 INPUT NODEFVAL data20
// Retrieval info: USED_PORT: data21 0 0 0 0 INPUT NODEFVAL data21
// Retrieval info: USED_PORT: data22 0 0 0 0 INPUT NODEFVAL data22
// Retrieval info: USED_PORT: data23 0 0 0 0 INPUT NODEFVAL data23
// Retrieval info: USED_PORT: data24 0 0 0 0 INPUT NODEFVAL data24
// Retrieval info: USED_PORT: data25 0 0 0 0 INPUT NODEFVAL data25
// Retrieval info: USED_PORT: data26 0 0 0 0 INPUT NODEFVAL data26
// Retrieval info: USED_PORT: data27 0 0 0 0 INPUT NODEFVAL data27
// Retrieval info: USED_PORT: data28 0 0 0 0 INPUT NODEFVAL data28
// Retrieval info: USED_PORT: data29 0 0 0 0 INPUT NODEFVAL data29
// Retrieval info: USED_PORT: data3 0 0 0 0 INPUT NODEFVAL data3
// Retrieval info: USED_PORT: data30 0 0 0 0 INPUT NODEFVAL data30
// Retrieval info: USED_PORT: data31 0 0 0 0 INPUT NODEFVAL data31
// Retrieval info: USED_PORT: data32 0 0 0 0 INPUT NODEFVAL data32
// Retrieval info: USED_PORT: data33 0 0 0 0 INPUT NODEFVAL data33
// Retrieval info: USED_PORT: data34 0 0 0 0 INPUT NODEFVAL data34
// Retrieval info: USED_PORT: data35 0 0 0 0 INPUT NODEFVAL data35
// Retrieval info: USED_PORT: data36 0 0 0 0 INPUT NODEFVAL data36
// Retrieval info: USED_PORT: data37 0 0 0 0 INPUT NODEFVAL data37
// Retrieval info: USED_PORT: data38 0 0 0 0 INPUT NODEFVAL data38
// Retrieval info: USED_PORT: data39 0 0 0 0 INPUT NODEFVAL data39
// Retrieval info: USED_PORT: data4 0 0 0 0 INPUT NODEFVAL data4
// Retrieval info: USED_PORT: data40 0 0 0 0 INPUT NODEFVAL data40
// Retrieval info: USED_PORT: data41 0 0 0 0 INPUT NODEFVAL data41
// Retrieval info: USED_PORT: data42 0 0 0 0 INPUT NODEFVAL data42
// Retrieval info: USED_PORT: data43 0 0 0 0 INPUT NODEFVAL data43
// Retrieval info: USED_PORT: data44 0 0 0 0 INPUT NODEFVAL data44
// Retrieval info: USED_PORT: data45 0 0 0 0 INPUT NODEFVAL data45
// Retrieval info: USED_PORT: data46 0 0 0 0 INPUT NODEFVAL data46
// Retrieval info: USED_PORT: data47 0 0 0 0 INPUT NODEFVAL data47
// Retrieval info: USED_PORT: data48 0 0 0 0 INPUT NODEFVAL data48
// Retrieval info: USED_PORT: data49 0 0 0 0 INPUT NODEFVAL data49
// Retrieval info: USED_PORT: data5 0 0 0 0 INPUT NODEFVAL data5
// Retrieval info: USED_PORT: data50 0 0 0 0 INPUT NODEFVAL data50
// Retrieval info: USED_PORT: data51 0 0 0 0 INPUT NODEFVAL data51
// Retrieval info: USED_PORT: data52 0 0 0 0 INPUT NODEFVAL data52
// Retrieval info: USED_PORT: data53 0 0 0 0 INPUT NODEFVAL data53
// Retrieval info: USED_PORT: data54 0 0 0 0 INPUT NODEFVAL data54
// Retrieval info: USED_PORT: data55 0 0 0 0 INPUT NODEFVAL data55
// Retrieval info: USED_PORT: data56 0 0 0 0 INPUT NODEFVAL data56
// Retrieval info: USED_PORT: data57 0 0 0 0 INPUT NODEFVAL data57
// Retrieval info: USED_PORT: data58 0 0 0 0 INPUT NODEFVAL data58
// Retrieval info: USED_PORT: data59 0 0 0 0 INPUT NODEFVAL data59
// Retrieval info: USED_PORT: data6 0 0 0 0 INPUT NODEFVAL data6
// Retrieval info: USED_PORT: data60 0 0 0 0 INPUT NODEFVAL data60
// Retrieval info: USED_PORT: data61 0 0 0 0 INPUT NODEFVAL data61
// Retrieval info: USED_PORT: data62 0 0 0 0 INPUT NODEFVAL data62
// Retrieval info: USED_PORT: data63 0 0 0 0 INPUT NODEFVAL data63
// Retrieval info: USED_PORT: data7 0 0 0 0 INPUT NODEFVAL data7
// Retrieval info: USED_PORT: data8 0 0 0 0 INPUT NODEFVAL data8
// Retrieval info: USED_PORT: data9 0 0 0 0 INPUT NODEFVAL data9
// Retrieval info: USED_PORT: result 0 0 0 0 OUTPUT NODEFVAL result
// Retrieval info: USED_PORT: sel 0 0 6 0 INPUT NODEFVAL sel[5..0]
// Retrieval info: CONNECT: result 0 0 0 0 @result 0 0 1 0
// Retrieval info: CONNECT: @data 0 0 1 63 data63 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 62 data62 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 61 data61 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 60 data60 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 59 data59 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 58 data58 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 57 data57 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 56 data56 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 55 data55 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 54 data54 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 53 data53 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 52 data52 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 51 data51 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 50 data50 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 49 data49 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 48 data48 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 47 data47 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 46 data46 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 45 data45 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 44 data44 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 43 data43 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 42 data42 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 41 data41 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 40 data40 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 39 data39 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 38 data38 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 37 data37 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 36 data36 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 35 data35 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 34 data34 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 33 data33 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 32 data32 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 31 data31 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 30 data30 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 29 data29 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 28 data28 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 27 data27 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 26 data26 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 25 data25 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 24 data24 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 23 data23 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 22 data22 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 21 data21 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 20 data20 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 19 data19 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 18 data18 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 17 data17 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 16 data16 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 15 data15 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 14 data14 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 13 data13 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 12 data12 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 11 data11 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 10 data10 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 9 data9 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 8 data8 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 7 data7 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 6 data6 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 5 data5 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 4 data4 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 3 data3 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 2 data2 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 1 data1 0 0 0 0
// Retrieval info: CONNECT: @data 0 0 1 0 data0 0 0 0 0
// Retrieval info: CONNECT: @sel 0 0 6 0 sel 0 0 6 0
// Retrieval info: LIBRARY: lpm lpm.lpm_components.all
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux641.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux641.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux641.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux641.bsf TRUE FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux641_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL lpm_mux641_bb.v TRUE
// Retrieval info: LIB_FILE: lpm
